
module adc_converter_IN2 (
	clk,
	reset_n,
	adc_data);	

	input		clk;
	input		reset_n;
	output	[11:0]	adc_data;
endmodule
