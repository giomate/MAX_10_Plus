// adc_converter_IN2.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module adc_converter_IN2 (
		output wire [11:0] adc_data, // adc_out.rx_in
		input  wire        clk,      //   clock.clk
		input  wire        reset_n   //   reset.reset_n
	);

	adc_converter_qip adc_in2_ch0_converter_0 (
		.clk      (clk),      //   clock.clk
		.reset_n  (reset_n),  //   reset.reset_n
		.adc_data (adc_data)  // adc_out.rx_in
	);

endmodule
