// anain2_converter.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module anain2_converter (
		input  wire        modular_adc_0_adc_pll_clock_clk,      //  modular_adc_0_adc_pll_clock.clk
		input  wire        modular_adc_0_adc_pll_locked_export,  // modular_adc_0_adc_pll_locked.export
		input  wire        modular_adc_0_clock_clk,              //          modular_adc_0_clock.clk
		input  wire        modular_adc_0_command_valid,          //        modular_adc_0_command.valid
		input  wire [4:0]  modular_adc_0_command_channel,        //                             .channel
		input  wire        modular_adc_0_command_startofpacket,  //                             .startofpacket
		input  wire        modular_adc_0_command_endofpacket,    //                             .endofpacket
		output wire        modular_adc_0_command_ready,          //                             .ready
		input  wire        modular_adc_0_reset_sink_reset_n,     //     modular_adc_0_reset_sink.reset_n
		output wire        modular_adc_0_response_valid,         //       modular_adc_0_response.valid
		output wire [4:0]  modular_adc_0_response_channel,       //                             .channel
		output wire [11:0] modular_adc_0_response_data,          //                             .data
		output wire        modular_adc_0_response_startofpacket, //                             .startofpacket
		output wire        modular_adc_0_response_endofpacket    //                             .endofpacket
	);

	anain2_converter_modular_adc_0 #(
		.is_this_first_or_second_adc (2)
	) modular_adc_0 (
		.clock_clk              (modular_adc_0_clock_clk),              //          clock.clk
		.reset_sink_reset_n     (modular_adc_0_reset_sink_reset_n),     //     reset_sink.reset_n
		.adc_pll_clock_clk      (modular_adc_0_adc_pll_clock_clk),      //  adc_pll_clock.clk
		.adc_pll_locked_export  (modular_adc_0_adc_pll_locked_export),  // adc_pll_locked.export
		.command_valid          (modular_adc_0_command_valid),          //        command.valid
		.command_channel        (modular_adc_0_command_channel),        //               .channel
		.command_startofpacket  (modular_adc_0_command_startofpacket),  //               .startofpacket
		.command_endofpacket    (modular_adc_0_command_endofpacket),    //               .endofpacket
		.command_ready          (modular_adc_0_command_ready),          //               .ready
		.response_valid         (modular_adc_0_response_valid),         //       response.valid
		.response_channel       (modular_adc_0_response_channel),       //               .channel
		.response_data          (modular_adc_0_response_data),          //               .data
		.response_startofpacket (modular_adc_0_response_startofpacket), //               .startofpacket
		.response_endofpacket   (modular_adc_0_response_endofpacket)    //               .endofpacket
	);

endmodule
