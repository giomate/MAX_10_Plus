
module adc_input2_channel0 (
	clk_clk,
	reset_reset_n,
	adc_in2_ch0_converter_0_adc_out_rx_in);	

	input		clk_clk;
	input		reset_reset_n;
	output	[11:0]	adc_in2_ch0_converter_0_adc_out_rx_in;
endmodule
