
module max_index_fft (
	clk_clk,
	reset_reset_n,
	index_fft_0_index_out_max_index_byte,
	index_fft_0_rx_input_rx_in);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	index_fft_0_index_out_max_index_byte;
	input	[11:0]	index_fft_0_rx_input_rx_in;
endmodule
