// tones_generator_sys.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module tones_generator_sys (
		input  wire        dac_tones_generator_0_clock_clk,            //    dac_tones_generator_0_clock.clk
		output wire [15:0] dac_tones_generator_0_dac_out_data_dac,     //  dac_tones_generator_0_dac_out.data_dac
		input  wire        dac_tones_generator_0_reset_reset_n,        //    dac_tones_generator_0_reset.reset_n
		output wire        dac_tones_generator_0_spi_data_data,        // dac_tones_generator_0_spi_data.data
		output wire        dac_tones_generator_0_spi_data_spi_clk,     //                               .spi_clk
		output wire        dac_tones_generator_0_spi_data_spi_sync,    //                               .spi_sync
		input  wire [4:0]  dac_tones_generator_0_switches_switches_in  // dac_tones_generator_0_switches.switches_in
	);

	tone_generator_qip dac_tones_generator_0 (
		.clk_in       (dac_tones_generator_0_clock_clk),            //    clock.clk
		.reset_n      (dac_tones_generator_0_reset_reset_n),        //    reset.reset_n
		.DAC_DATA     (dac_tones_generator_0_spi_data_data),        // spi_data.data
		.DAC_SCLK     (dac_tones_generator_0_spi_data_spi_clk),     //         .spi_clk
		.DAC_SYNC_n   (dac_tones_generator_0_spi_data_spi_sync),    //         .spi_sync
		.SW           (dac_tones_generator_0_switches_switches_in), // switches.switches_in
		.dac_data_out (dac_tones_generator_0_dac_out_data_dac)      //  dac_out.data_dac
	);

endmodule
