
module fft_loop_test (
	clk_clk,
	index_fft_0_index_out_max_index_byte,
	pio_0_external_connection_export,
	reset_reset_n,
	dac_tones_generator_0_spi_data_data,
	dac_tones_generator_0_spi_data_spi_clk,
	dac_tones_generator_0_spi_data_spi_sync,
	dac_tones_generator_0_switches_switches_in);	

	input		clk_clk;
	output	[7:0]	index_fft_0_index_out_max_index_byte;
	output	[7:0]	pio_0_external_connection_export;
	input		reset_reset_n;
	output		dac_tones_generator_0_spi_data_data;
	output		dac_tones_generator_0_spi_data_spi_clk;
	output		dac_tones_generator_0_spi_data_spi_sync;
	input	[4:0]	dac_tones_generator_0_switches_switches_in;
endmodule
